*** SPICE deck for cell INV{lay} from library InverterProject
*** Created on Fri May 10, 2024 13:23:57
*** Last revised on Mon May 27, 2024 12:59:43
*** Written on Mon May 27, 2024 12:59:51 by Electric VLSI Design System, version 9.07
*** Layout tech: mocmos, foundry MOSIS
*** UC SPICE *** , MIN_RESIST 4.0, MIN_CAPAC 0.1FF

*** TOP LEVEL CELL: InverterProject:INV{lay}
Mnmos@0 gnd in out gnd NMOS L=1.2U W=6U AS=46.44P AD=84.24P PS=45.6U PD=74.4U
Mpmos@0 vdd in out vdd PMOS L=1.2U W=12U AS=46.44P AD=113.04P PS=45.6U PD=98.4U

* Spice Code nodes in cell cell 'InverterProject:INV{lay}'
vdd vdd 0 DC 5
vin in 0 pwl 5n 0 10n 0 20n 5 50n 5 60n 0 70n 0 80n 0 100n 0
cload out 0 250fF
.measure tran tf trig v(out) val= 4.5 fall=1 td=1ns targ v(out) val=0.5 fall=1
.measure tran tr trig v(out) val= 0.5 rise=1 td=5ns targ v(out) val=4.5 rise=1
.tran 0 0.1us
.include C:\LTspice\C5_models.txt
.END
